module MIPS #(
    parameters
) (
    ports
);
    
endmodule