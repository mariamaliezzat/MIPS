module Register_File (
                       input [31:0] WD3,
                       input [4:0] A1,
                       input [4:0] A2,
                       input [4:0] A3,
                       input reset_b,
                       input clk,
                       output [31:0] RD1,
                       output [31:0] RD2
);

reg [31:0] register_file [99:0];
reg WE3;
integer i; 
always@(posedge clk)

begin
if(reset_b)
begin
if(WD3==1)
register_file[A3] <= WD3;
end
else
begin
for(i=0;i<32;i=i+1)
begin
register_file[i] <=0;
end
end

end


assign RD1=register_file[A1];
assign RD2=register_file[A2];




endmodule